module xor4 ();
p


endmodule:
